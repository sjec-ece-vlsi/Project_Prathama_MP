/*
 RAM has 16K memory loaction with 16 bit width. 
 Use parameter to define Location, width and address bits required for the ROM.
*/

module RAM_16k(
  
);
  
// parameter for Address width, Data_bus and Memeory Depth or locations
  
// Declare inputs and outputs including control signals
  
  
// Declare Required internal wires or registers
  
  
 // Logic goes here
  
  
  //end of the logic
  
  
endmodule
