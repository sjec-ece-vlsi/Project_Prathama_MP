/*
 Create  a testbench to test 8k ROM with Control signals
 

*/
module rom_tb();
  
  // Declare required registers, wires and parameters for Device under test (DUT) 
  
  // Call for DUT
  
  
  // Initial blocks
  
  
  //
  
  // Verfication code 
  
  
  //
  
  //end of logic
  
endmodule
