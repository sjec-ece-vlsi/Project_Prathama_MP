/*
 Create  a testbench to test 16k RAM with Control signals
 
*/
module RAM_tb();
  
  // Declare required registers, wires and parameters for Device under test (DUT) 
  
  // Call for DUT
  
  
  // Initial blocks
  
  
  //
  
  // Verfication code 
  
  
  //
  
  //end of logic
  
endmodule
