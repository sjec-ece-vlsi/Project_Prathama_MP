module ROM_8k(
  input cs
