module RAM_16k(
  
