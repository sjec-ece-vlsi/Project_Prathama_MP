module ROM_8k(
  
);
  
  
  
endmodule
